AOI
Vdd	vdd	0	5
VinA nga	0 PULSE( 5, 0, 0, 1u, 1u, 4.998m, 10m )
VinB ngb	0 PULSE( 5, 0, 0, 1u, 1u, 2.5m, 5m )
VinBi ngbi	0 PULSE( 0, 5, 0, 1u, 1u, 2.5m, 5m ); supplies
VinC ngc	0 PULSE( 5, 0, 0, 1u, 1u, 1.248m, 2.5m )
VinD ngd	0 PULSE( 5, 0, 0, 1u, 1u, 0.627m, 1.25m )

*std width = 4u std N length = 7.8u	std P length =2u
MAP		vdd		nga		ND		vdd		MP	W=2u		L=1u
MBPI	vdd		ngbi	ndCP	vdd		MP	W=2u		L=0.5u
MCP		ndCP	ngc		ND		vdd		MP	W=2u		L=0.5u; PMOS
MDP		ND		ngd		ndout	vdd		MP	W=2u		L=1u
MBP		ND		ngb		ndout	vdd		MP	W=2u		L=1u

MAN		ndout	nga		ndbic	0		MN	W=2u		L=3.9u
MBIN	ndbic	ngbi	0		0		MN	W=1u		L=3.9u
MCN		ndbic	ngc		0		0		MN	W=1u		L=3.9u;NMOS
MDN		ndout	ngd		ndbn	0		MN	W=2u		L=3.9u
MBN		ndbn	ngb		0		0		MN	W=2u		L=3.9u

*inverter
MPin	vdd		ndout	out		vdd	MP	W=4u	L=2u
MNin	out		ndout	0		0	MN	W=4u	L=7.8u


.lib tsmc035.lib
.tran	1e-03	0.1e-1
.end
